// i2c_controller_avmm_bridge.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module i2c_controller_avmm_bridge (
		input  wire        i2c_clock_clk,     //  i2c_clock.clk
		input  wire [3:0]  i2c_csr_address,   //    i2c_csr.address
		input  wire        i2c_csr_read,      //           .read
		input  wire        i2c_csr_write,     //           .write
		input  wire [31:0] i2c_csr_writedata, //           .writedata
		output wire [31:0] i2c_csr_readdata,  //           .readdata
		output wire        i2c_irq_irq,       //    i2c_irq.irq
		input  wire        i2c_reset_reset_n, //  i2c_reset.reset_n
		input  wire        i2c_serial_sda_in, // i2c_serial.sda_in
		input  wire        i2c_serial_scl_in, //           .scl_in
		output wire        i2c_serial_sda_oe, //           .sda_oe
		output wire        i2c_serial_scl_oe  //           .scl_oe
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (64),
		.FIFO_DEPTH_LOG2 (6)
	) i2c_master (
		.clk       (i2c_clock_clk),        //            clock.clk
		.rst_n     (i2c_reset_reset_n),    //       reset_sink.reset_n
		.intr      (i2c_irq_irq),          // interrupt_sender.irq
		.addr      (i2c_csr_address),      //              csr.address
		.read      (i2c_csr_read),         //                 .read
		.write     (i2c_csr_write),        //                 .write
		.writedata (i2c_csr_writedata),    //                 .writedata
		.readdata  (i2c_csr_readdata),     //                 .readdata
		.sda_in    (i2c_serial_sda_in),    //       i2c_serial.sda_in
		.scl_in    (i2c_serial_scl_in),    //                 .scl_in
		.sda_oe    (i2c_serial_sda_oe),    //                 .sda_oe
		.scl_oe    (i2c_serial_scl_oe),    //                 .scl_oe
		.src_data  (),                     //      (terminated)
		.src_valid (),                     //      (terminated)
		.src_ready (1'b0),                 //      (terminated)
		.snk_data  (16'b0000000000000000), //      (terminated)
		.snk_valid (1'b0),                 //      (terminated)
		.snk_ready ()                      //      (terminated)
	);

endmodule
