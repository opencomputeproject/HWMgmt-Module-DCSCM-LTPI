
package ltpi_data_channel_controller_model_pkg;
    `include "ltpi_data_channel_controller_driver.svh"
endpackage
