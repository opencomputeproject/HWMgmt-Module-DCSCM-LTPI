
package I2C_controller_bridge_pkg;
    `include "I2C_controller_bridge_driver.svh"
endpackage
